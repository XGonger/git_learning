module tb;
  wire a;
  wire b;

endmodule
